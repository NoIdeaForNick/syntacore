module cross_bar(  
                    

);